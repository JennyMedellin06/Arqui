library verilog;
use verilog.vl_types.all;
entity Control is
    port(
        OP              : in     vl_logic_vector(5 downto 0);
        RegDst          : out    vl_logic;
        BranchEQ        : out    vl_logic;
        BranchNE        : out    vl_logic;
        MemRead         : out    vl_logic;
        MemtoReg        : out    vl_logic;
        MemWrite        : out    vl_logic;
        ALUSrc          : out    vl_logic;
        RegWrite        : out    vl_logic;
        ALUOp           : out    vl_logic_vector(3 downto 0)
    );
end Control;
